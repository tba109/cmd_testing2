library verilog;
use verilog.vl_types.all;
entity phf_testing_tb is
end phf_testing_tb;
