library verilog;
use verilog.vl_types.all;
entity cmd_testing2_tb is
end cmd_testing2_tb;
