`ifndef _CMD_DEFS_VH_
`define _CMD_DEFS_VH_

`define N_TAP_CTL_SIZE 18

`endif
